`timescale 1ns/1ns

// FIFO Parameters 
`define     FIFO_WIDTH          8
`define     FIFO_DEPTH          16
`define     FIFO_ADDR_WIDTH     (1+4)   // one for MSB 