`include "defines.vh"

module FIFOSync (
    input wire clk,
    input wire restn,
    input wire [`FIFO_ADDR_WIDTH-1: 0] ptr_in,
    output wire [`FIFO_ADDR_WIDTH-1: 0] ptr_out
);



endmodule